test markus
