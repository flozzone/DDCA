test markus
test florin
test2 markus
