test markus
test florin
