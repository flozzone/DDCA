test markus
test florin
test2 markus
test3 markus
-------------
florin
petar
