1337hetti
