1337hetti
added line